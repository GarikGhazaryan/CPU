module Ham ()

wire [3:0] in_dat
wire [i6:0] ham_dat;




encod en (data_in, data_h_out);

decod de (data_h_in, data_out);
